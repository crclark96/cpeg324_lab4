-------------------------------------------------------------------------------
-- Title      : comparator_2_bit
-- Project    : 
-------------------------------------------------------------------------------
-- File       : comparator_2_bit.vhdl
-- Author     : Collin Clark  <collinclark@wifi-roaming-128-4-61-116.host.udel.edu>
-- Company    : 
-- Created    : 2018-05-12
-- Last update: 2018-05-12
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2018 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2018-05-12  1.0      collinclark     Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------

entity comparator_2_bit is

  port (a     : in  std_logic_vector(1 downto 0);
        b     : in  std_logic_vector(1 downto 0);
        s     : out std_logic
        );

end entity comparator_2_bit;

-------------------------------------------------------------------------------

architecture str of comparator_2_bit is

  -----------------------------------------------------------------------------
  -- Internal signal declarations
  -----------------------------------------------------------------------------

begin  -- architecture str

  -----------------------------------------------------------------------------
  -- Component instantiations
  -----------------------------------------------------------------------------

  s <= not ((a(0) xor b(0)) or (a(1) xor b(1)));
  
  
end architecture str;

-------------------------------------------------------------------------------
